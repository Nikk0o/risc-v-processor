`ifndef ALUOP_H
`define ALUOP_H

`define NONE 0
`define ADD 1
`define SUB 2
`define AND 3
`define XOR 4
`define XNOR 5
`define OR 6
`define NOT 7
`define LSHIFT 8
`define ARSHIFT 9
`define LRSHIFT 10
`define MUL 11
`define DIV 12
`define SUBU 13
`define DIVU 14
`define REMU 15

`endif
